* SPICE3 file created from 41osu.ext - technology: scmos

.option scale=0.1u

.include NMOS-180nm.lib
.include PMOS-180nm.lib

M1000 a_26_n68# S0 I3 vss nfet w=8 l=2
+  ad=184 pd=94 as=56 ps=30
M1001 a_26_69# S0bar I0 vss nfet w=8 l=2
+  ad=184 pd=94 as=56 ps=30
M1002 outpt S1 a_26_n68# vss nfet w=8 l=2
+  ad=128 pd=64 as=0 ps=0
M1003 vcc S0 S0bar w_n32_136# pfet w=8 l=2
+  ad=168 pd=90 as=64 ps=32
M1004 a_26_69# S0bar I1 w_11_91# pfet w=8 l=2
+  ad=184 pd=94 as=56 ps=30
M1005 a_96_n20# S1 vss vss nfet w=8 l=2
+  ad=64 pd=32 as=168 ps=90
M1006 a_26_n68# a_n26_n20# I3 w_11_n46# pfet w=8 l=2
+  ad=184 pd=94 as=56 ps=30
M1007 outpt a_96_n20# a_26_n68# w_133_n46# pfet w=8 l=2
+  ad=128 pd=64 as=0 ps=0
M1008 a_26_69# S0 I0 w_11_145# pfet w=8 l=2
+  ad=0 pd=0 as=56 ps=30
M1009 vcc S0 a_n26_n20# w_n32_n1# pfet w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1010 a_26_n68# S0 I2 w_11_8# pfet w=8 l=2
+  ad=0 pd=0 as=56 ps=30
M1011 a_26_n68# a_n26_n20# I2 vss nfet w=8 l=2
+  ad=0 pd=0 as=56 ps=30
M1012 outpt a_96_n20# a_26_69# vss nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 outpt S1 a_26_69# w_133_8# pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 S0bar S0 vss vss nfet w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1015 a_n26_n20# S0 vss vss nfet w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1016 vcc S1 a_96_n20# w_90_n1# pfet w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1017 a_26_69# S0 I1 vss nfet w=8 l=2
+  ad=0 pd=0 as=56 ps=30
C0 S0 vss 3.93fF


V1 vcc 0 .5
V2 S0 0 PULSE(.5 -.5 0.1n 0.1n 0.1n 2u 4u)
V3 S1 0 PULSE(.5 -.5 0.1n 0.1n 0.1n 4u 8u)
V4 I0 0 1.235
V5 I1 0 PULSE(1 .5 0.1n 0.1n 0.1n 0.8u 1.6u)
V6 I2 0 1.235
V7 I3 0 PULSE(1 .5 0.1n 0.1n 0.1n 0.8u 1.6u)
V8 vss 0 -0.5
.tran 0.001u 10u
.control
run
plot V(S0)
plot V(S1)
plot V(I0)
plot V(I1)
plot V(I2)
plot V(I3)
plot V(outpt)
plot V(S0bar)
.endc
.end41

* SPICE3 file created from 21try.ext - technology: scmos

.option scale=0.1u
.include NMOS-180nm.lib
.include PMOS-180nm.lib

M1000 out a_n42_n33# I0 vss nfet w=14 l=2
+  ad=392 pd=112 as=196 ps=56
M1001 out sel I1 vss nfet w=14 l=2
+  ad=0 pd=0 as=196 ps=56
M1002 a_n42_n33# sel vcc w_n62_5# pfet w=14 l=2
+  ad=182 pd=54 as=210 ps=58
M1003 out a_n42_n33# I1 w_n62_5# pfet w=14 l=2
+  ad=392 pd=112 as=196 ps=56
M1004 out sel I0 w_n62_5# pfet w=14 l=2
+  ad=0 pd=0 as=196 ps=56
M1005 a_n42_n33# sel vss vss nfet w=14 l=2
+  ad=182 pd=54 as=210 ps=58
C0 w_n62_5# vss 2.64fF

V1 vcc 0 1
V2 sel 0 PULSE(.5 -.5 0.1n 0.1n 0.1n 10u 20u)
V4 I0 0 SINE(0 1 800000)	
V5 I1 0 2.5
V8 vss 0 -1
.tran 0.001u 30u
.control
run
plot V(sel)
plot V(I0)
plot V(I1)
plot V(out)
.endc
.end

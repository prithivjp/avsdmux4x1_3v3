magic
tech scmos
timestamp 1594202356
<< nwell >>
rect 9 25 91 45
rect -18 -1 104 19
<< ntransistor >>
rect 22 52 24 60
rect 41 52 43 60
rect 76 52 78 60
rect -3 -16 -1 -8
rect 16 -16 18 -8
rect 41 -16 43 -8
rect 66 -16 68 -8
rect 85 -16 87 -8
<< ptransistor >>
rect 22 31 24 39
rect 41 31 43 39
rect 76 31 78 39
rect -3 5 -1 13
rect 16 5 18 13
rect 41 5 43 13
rect 66 5 68 13
rect 85 5 87 13
<< ndiffusion >>
rect 15 58 22 60
rect 15 54 17 58
rect 21 54 22 58
rect 15 52 22 54
rect 24 58 31 60
rect 24 54 25 58
rect 29 54 31 58
rect 24 52 31 54
rect 34 59 41 60
rect 34 55 36 59
rect 40 55 41 59
rect 34 52 41 55
rect 43 58 50 60
rect 43 54 44 58
rect 48 54 50 58
rect 43 52 50 54
rect 69 58 76 60
rect 69 54 71 58
rect 75 54 76 58
rect 69 52 76 54
rect 78 58 85 60
rect 78 54 79 58
rect 83 54 85 58
rect 78 52 85 54
rect -10 -10 -3 -8
rect -10 -14 -8 -10
rect -4 -14 -3 -10
rect -10 -16 -3 -14
rect -1 -10 6 -8
rect -1 -14 0 -10
rect 4 -14 6 -10
rect -1 -16 6 -14
rect 9 -10 16 -8
rect 9 -14 11 -10
rect 15 -14 16 -10
rect 9 -16 16 -14
rect 18 -10 25 -8
rect 18 -14 19 -10
rect 23 -14 25 -10
rect 18 -16 25 -14
rect 34 -11 41 -8
rect 34 -15 36 -11
rect 40 -15 41 -11
rect 34 -16 41 -15
rect 43 -10 50 -8
rect 43 -14 44 -10
rect 48 -14 50 -10
rect 43 -16 50 -14
rect 59 -10 66 -8
rect 59 -14 61 -10
rect 65 -14 66 -10
rect 59 -16 66 -14
rect 68 -10 75 -8
rect 68 -14 69 -10
rect 73 -14 75 -10
rect 68 -16 75 -14
rect 78 -10 85 -8
rect 78 -14 80 -10
rect 84 -14 85 -10
rect 78 -16 85 -14
rect 87 -10 94 -8
rect 87 -14 88 -10
rect 92 -14 94 -10
rect 87 -16 94 -14
<< pdiffusion >>
rect 15 37 22 39
rect 15 33 17 37
rect 21 33 22 37
rect 15 31 22 33
rect 24 37 31 39
rect 24 33 25 37
rect 29 33 31 37
rect 24 31 31 33
rect 34 36 41 39
rect 34 32 36 36
rect 40 32 41 36
rect 34 31 41 32
rect 43 37 50 39
rect 43 33 44 37
rect 48 33 50 37
rect 43 31 50 33
rect 69 37 76 39
rect 69 33 71 37
rect 75 33 76 37
rect 69 31 76 33
rect 78 37 85 39
rect 78 33 79 37
rect 83 33 85 37
rect 78 31 85 33
rect -10 11 -3 13
rect -10 7 -8 11
rect -4 7 -3 11
rect -10 5 -3 7
rect -1 11 6 13
rect -1 7 0 11
rect 4 7 6 11
rect -1 5 6 7
rect 9 11 16 13
rect 9 7 11 11
rect 15 7 16 11
rect 9 5 16 7
rect 18 11 25 13
rect 18 7 19 11
rect 23 7 25 11
rect 18 5 25 7
rect 34 12 41 13
rect 34 8 36 12
rect 40 8 41 12
rect 34 5 41 8
rect 43 11 50 13
rect 43 7 44 11
rect 48 7 50 11
rect 43 5 50 7
rect 59 11 66 13
rect 59 7 61 11
rect 65 7 66 11
rect 59 5 66 7
rect 68 11 75 13
rect 68 7 69 11
rect 73 7 75 11
rect 68 5 75 7
rect 78 11 85 13
rect 78 7 80 11
rect 84 7 85 11
rect 78 5 85 7
rect 87 11 94 13
rect 87 7 88 11
rect 92 7 94 11
rect 87 5 94 7
<< ndcontact >>
rect 17 54 21 58
rect 25 54 29 58
rect 36 55 40 59
rect 44 54 48 58
rect 71 54 75 58
rect 79 54 83 58
rect -8 -14 -4 -10
rect 0 -14 4 -10
rect 11 -14 15 -10
rect 19 -14 23 -10
rect 36 -15 40 -11
rect 44 -14 48 -10
rect 61 -14 65 -10
rect 69 -14 73 -10
rect 80 -14 84 -10
rect 88 -14 92 -10
<< pdcontact >>
rect 17 33 21 37
rect 25 33 29 37
rect 36 32 40 36
rect 44 33 48 37
rect 71 33 75 37
rect 79 33 83 37
rect -8 7 -4 11
rect 0 7 4 11
rect 11 7 15 11
rect 19 7 23 11
rect 36 8 40 12
rect 44 7 48 11
rect 61 7 65 11
rect 69 7 73 11
rect 80 7 84 11
rect 88 7 92 11
<< psubstratepcontact >>
rect 36 64 40 68
rect 36 -29 40 -25
<< nsubstratencontact >>
rect 36 20 40 24
<< polysilicon >>
rect 22 60 24 63
rect 41 62 78 64
rect 41 60 43 62
rect 76 60 78 62
rect 22 51 24 52
rect 22 49 34 51
rect 22 39 24 42
rect 41 39 43 52
rect 50 48 72 50
rect 76 49 78 52
rect 70 44 72 48
rect 70 42 78 44
rect 76 39 78 42
rect 22 30 24 31
rect 41 30 43 31
rect 22 28 43 30
rect 76 28 78 31
rect 41 27 43 28
rect -3 13 -1 17
rect 16 15 68 17
rect 16 13 18 15
rect 41 13 43 15
rect 66 13 68 15
rect 85 13 87 17
rect -3 -1 -1 5
rect -3 -3 8 -1
rect 16 -2 18 5
rect 6 -5 8 -3
rect 26 -5 32 -3
rect -3 -8 -1 -6
rect 6 -7 28 -5
rect 16 -8 18 -7
rect 41 -8 43 5
rect 66 -2 68 5
rect 85 -1 87 5
rect 77 -3 87 -1
rect 52 -5 60 -3
rect 77 -5 79 -3
rect 58 -7 79 -5
rect 66 -8 68 -7
rect 85 -8 87 -6
rect -3 -22 -1 -16
rect 16 -18 18 -16
rect 41 -22 43 -16
rect 66 -18 68 -16
rect 85 -22 87 -16
rect -3 -24 87 -22
<< polycontact >>
rect 34 47 38 51
rect 46 47 50 51
rect 32 -6 36 -2
rect 48 -6 52 -2
<< metal1 >>
rect -23 -29 -19 75
rect 25 71 75 75
rect 25 58 29 71
rect 17 49 21 54
rect 3 45 21 49
rect 3 24 7 45
rect 17 37 21 45
rect 40 65 58 68
rect 36 59 40 64
rect 25 37 29 54
rect 44 51 48 54
rect 38 47 46 51
rect 44 37 48 47
rect 36 24 40 32
rect 0 20 15 24
rect 0 11 4 20
rect -8 -10 -4 7
rect 0 -10 4 7
rect 11 11 15 20
rect 26 20 36 24
rect 40 20 44 24
rect 11 -10 15 7
rect 19 -10 23 7
rect 26 -29 29 20
rect 36 12 40 20
rect 44 -2 48 7
rect 36 -6 48 -2
rect 44 -10 48 -6
rect -23 -33 29 -29
rect 36 -25 40 -15
rect 55 -29 58 65
rect 71 58 75 71
rect 71 37 75 54
rect 79 49 83 54
rect 79 45 97 49
rect 79 37 83 45
rect 93 24 97 45
rect 69 20 97 24
rect 69 11 73 20
rect 61 -10 65 7
rect 69 -10 73 7
rect 80 11 84 20
rect 80 -10 84 7
rect 88 -10 92 7
rect 105 -29 109 75
rect 36 -33 109 -29
rect -23 -37 -19 -33
rect 105 -37 109 -33
<< labels >>
rlabel metal1 21 -3 21 -3 1 I0
rlabel metal1 -6 -4 -6 -4 1 I1
rlabel metal1 63 -3 63 -3 1 I2
rlabel metal1 90 -4 90 -4 1 I3
rlabel polysilicon 42 46 42 46 1 S1
rlabel polysilicon 42 -7 42 -7 1 S0
rlabel metal1 50 73 50 73 5 out
rlabel metal1 107 22 107 22 7 VSS
rlabel metal1 -21 24 -21 24 3 VDD
<< end >>

* C:\Users\prith\Desktop\check\Data Acquisition System.asc
M1 I0 sbar N001 vee n_mos l=0.18u w=0.36u
M2 I1 S0 N001 vee n_mos l=0.18u w=0.36u
M3 N001 S0 I0 vdd p_mos l=0.18u w=0.9u
M4 N001 sbar I1 vdd p_mos l=0.18u w=0.9u
M5 vcc S0 sbar vdd p_mos l=0.18u w=0.9u
M6 sbar S0 vss vee n_mos l=0.18u w=0.36u
V1 vdd 0 1.6
V2 vee 0 -1
V3 vcc 0 1
V4 vss 0 -1
V5 S0 0 PULSE(.5 -.5 0.1n 0.1n 0.1n 1u 2u)
V6 I0 0 SINE(0 1 25000000)
V7 I1 0 .5
M11 N001 N002 outpt vee n_mos l=0.18u w=0.36u
M12 N003 S1 outpt vee n_mos l=0.18u w=0.36u
M13 outpt S1 N001 vdd p_mos l=0.18u w=0.9u
M14 outpt N002 N003 vdd p_mos l=0.18u w=0.9u
M15 vcc S1 N002 vdd p_mos l=0.18u w=0.9u
M16 N002 S1 vss vee n_mos l=0.18u w=0.36u
M17 I2 sbar N003 vee n_mos l=0.18u w=0.36u
M18 I3 S0 N003 vee n_mos l=0.18u w=0.36u
M19 N003 S0 I2 vdd p_mos l=0.18u w=0.9u
M20 N003 sbar I3 vdd p_mos l=0.18u w=0.9u
V9 I3 0 .7
V10 S1 0 PULSE(.5 -.5 0.1n 0.1n 0.1n 2u 4u)
V11 I2 0 PULSE(-1 1 0.0001n 0.0001n 0.0001n 0.1u 0.2u)
.model NMOS NMOS
.model PMOS PMOS

.tran 0.001u 4u
.inc osulib.lib
.control
run
plot v(outpt)
.endc
.end

magic
tech scmos
timestamp 1593430242
<< nwell >>
rect -32 136 -12 165
rect 11 145 40 165
rect 11 91 40 111
rect -32 -1 -12 28
rect 11 8 40 28
rect 90 -1 110 28
rect 133 8 162 28
rect 11 -46 40 -26
rect 133 -46 162 -26
<< ntransistor >>
rect 24 123 26 131
rect -26 115 -18 117
rect 24 69 26 77
rect 24 -14 26 -6
rect -26 -22 -18 -20
rect 146 -14 148 -6
rect 96 -22 104 -20
rect 24 -68 26 -60
rect 146 -68 148 -60
<< ptransistor >>
rect -26 150 -18 152
rect 24 151 26 159
rect 24 97 26 105
rect -26 13 -18 15
rect 24 14 26 22
rect 96 13 104 15
rect 146 14 148 22
rect 24 -40 26 -32
rect 146 -40 148 -32
<< ndiffusion >>
rect -26 124 -18 125
rect -26 120 -24 124
rect -20 120 -18 124
rect -26 117 -18 120
rect 17 129 24 131
rect 17 124 18 129
rect 23 124 24 129
rect 17 123 24 124
rect 26 129 34 131
rect 26 124 27 129
rect 32 124 34 129
rect 26 123 34 124
rect -26 113 -18 115
rect -26 109 -24 113
rect -20 109 -18 113
rect -26 108 -18 109
rect 17 75 24 77
rect 17 70 18 75
rect 23 70 24 75
rect 17 69 24 70
rect 26 75 34 77
rect 26 70 27 75
rect 32 70 34 75
rect 26 69 34 70
rect -26 -13 -18 -12
rect -26 -17 -24 -13
rect -20 -17 -18 -13
rect -26 -20 -18 -17
rect 17 -8 24 -6
rect 17 -13 18 -8
rect 23 -13 24 -8
rect 17 -14 24 -13
rect 26 -8 34 -6
rect 26 -13 27 -8
rect 32 -13 34 -8
rect 26 -14 34 -13
rect -26 -24 -18 -22
rect -26 -28 -24 -24
rect -20 -28 -18 -24
rect -26 -29 -18 -28
rect 96 -13 104 -12
rect 96 -17 98 -13
rect 102 -17 104 -13
rect 96 -20 104 -17
rect 139 -8 146 -6
rect 139 -13 140 -8
rect 145 -13 146 -8
rect 139 -14 146 -13
rect 148 -8 156 -6
rect 148 -13 149 -8
rect 154 -13 156 -8
rect 148 -14 156 -13
rect 96 -24 104 -22
rect 96 -28 98 -24
rect 102 -28 104 -24
rect 96 -29 104 -28
rect 17 -62 24 -60
rect 17 -67 18 -62
rect 23 -67 24 -62
rect 17 -68 24 -67
rect 26 -62 34 -60
rect 26 -67 27 -62
rect 32 -67 34 -62
rect 26 -68 34 -67
rect 139 -62 146 -60
rect 139 -67 140 -62
rect 145 -67 146 -62
rect 139 -68 146 -67
rect 148 -62 156 -60
rect 148 -67 149 -62
rect 154 -67 156 -62
rect 148 -68 156 -67
<< pdiffusion >>
rect -26 158 -18 159
rect -26 154 -24 158
rect -20 154 -18 158
rect -26 152 -18 154
rect 17 157 24 159
rect 17 152 18 157
rect 23 152 24 157
rect 17 151 24 152
rect 26 157 34 159
rect 26 152 27 157
rect 32 152 34 157
rect 26 151 34 152
rect -26 147 -18 150
rect -26 143 -24 147
rect -20 143 -18 147
rect -26 142 -18 143
rect 17 103 24 105
rect 17 98 18 103
rect 23 98 24 103
rect 17 97 24 98
rect 26 103 34 105
rect 26 98 27 103
rect 32 98 34 103
rect 26 97 34 98
rect -26 21 -18 22
rect -26 17 -24 21
rect -20 17 -18 21
rect -26 15 -18 17
rect 17 20 24 22
rect 17 15 18 20
rect 23 15 24 20
rect 17 14 24 15
rect 26 20 34 22
rect 26 15 27 20
rect 32 15 34 20
rect 96 21 104 22
rect 96 17 98 21
rect 102 17 104 21
rect 96 15 104 17
rect 26 14 34 15
rect -26 10 -18 13
rect -26 6 -24 10
rect -20 6 -18 10
rect -26 5 -18 6
rect 139 20 146 22
rect 139 15 140 20
rect 145 15 146 20
rect 139 14 146 15
rect 148 20 156 22
rect 148 15 149 20
rect 154 15 156 20
rect 148 14 156 15
rect 96 10 104 13
rect 96 6 98 10
rect 102 6 104 10
rect 96 5 104 6
rect 17 -34 24 -32
rect 17 -39 18 -34
rect 23 -39 24 -34
rect 17 -40 24 -39
rect 26 -34 34 -32
rect 26 -39 27 -34
rect 32 -39 34 -34
rect 26 -40 34 -39
rect 139 -34 146 -32
rect 139 -39 140 -34
rect 145 -39 146 -34
rect 139 -40 146 -39
rect 148 -34 156 -32
rect 148 -39 149 -34
rect 154 -39 156 -34
rect 148 -40 156 -39
<< ndcontact >>
rect -24 120 -20 124
rect 18 124 23 129
rect 27 124 32 129
rect -24 109 -20 113
rect 18 70 23 75
rect 27 70 32 75
rect -24 -17 -20 -13
rect 18 -13 23 -8
rect 27 -13 32 -8
rect -24 -28 -20 -24
rect 98 -17 102 -13
rect 140 -13 145 -8
rect 149 -13 154 -8
rect 98 -28 102 -24
rect 18 -67 23 -62
rect 27 -67 32 -62
rect 140 -67 145 -62
rect 149 -67 154 -62
<< pdcontact >>
rect -24 154 -20 158
rect 18 152 23 157
rect 27 152 32 157
rect -24 143 -20 147
rect 18 98 23 103
rect 27 98 32 103
rect -24 17 -20 21
rect 18 15 23 20
rect 27 15 32 20
rect 98 17 102 21
rect -24 6 -20 10
rect 140 15 145 20
rect 149 15 154 20
rect 98 6 102 10
rect 18 -39 23 -34
rect 27 -39 32 -34
rect 140 -39 145 -34
rect 149 -39 154 -34
<< psubstratepcontact >>
rect -30 93 -26 97
rect -18 93 -14 97
rect -30 -44 -26 -40
rect -18 -44 -14 -40
rect 92 -44 96 -40
rect 104 -44 108 -40
<< nsubstratencontact >>
rect -30 170 -26 174
rect -18 170 -14 174
rect -30 33 -26 37
rect -18 33 -14 37
rect 92 33 96 37
rect 104 33 108 37
<< polysilicon >>
rect 2 168 26 170
rect 2 152 4 168
rect 24 159 26 168
rect -38 150 -26 152
rect -18 150 4 152
rect -38 136 -36 150
rect 24 142 26 151
rect -44 134 -36 136
rect -44 56 -42 134
rect -38 117 -36 134
rect -6 128 2 132
rect 24 131 26 134
rect 0 118 2 128
rect 24 118 26 123
rect -38 115 -26 117
rect -18 115 -6 117
rect 0 116 26 118
rect -8 112 -6 115
rect -8 110 4 112
rect 2 66 4 110
rect 24 105 26 116
rect 24 88 26 97
rect 24 77 26 80
rect 24 66 26 69
rect 2 64 26 66
rect -50 54 -42 56
rect -44 -4 -42 54
rect 2 31 26 33
rect 2 15 4 31
rect 24 22 26 31
rect 124 31 148 33
rect -38 13 -26 15
rect -18 13 4 15
rect 124 15 126 31
rect 146 22 148 31
rect -38 -4 -36 13
rect 24 5 26 14
rect 84 13 96 15
rect 104 13 126 15
rect 84 -2 86 13
rect 146 5 148 14
rect -44 -6 -36 -4
rect -38 -20 -36 -6
rect -6 -9 2 -5
rect 24 -6 26 -3
rect 78 -4 86 -2
rect 0 -19 2 -9
rect 24 -19 26 -14
rect -38 -22 -26 -20
rect -18 -22 -6 -20
rect 0 -21 26 -19
rect -8 -25 -6 -22
rect -8 -27 4 -25
rect 2 -71 4 -27
rect 24 -32 26 -21
rect 84 -20 86 -4
rect 116 -9 124 -5
rect 146 -6 148 -3
rect 122 -19 124 -9
rect 146 -19 148 -14
rect 84 -22 96 -20
rect 104 -22 116 -20
rect 122 -21 148 -19
rect 114 -25 116 -22
rect 114 -27 126 -25
rect 24 -49 26 -40
rect 24 -60 26 -57
rect 24 -71 26 -68
rect 2 -73 26 -71
rect 124 -71 126 -27
rect 146 -32 148 -21
rect 146 -49 148 -40
rect 146 -60 148 -57
rect 146 -71 148 -68
rect 124 -73 148 -71
<< polycontact >>
rect -10 128 -6 132
rect -10 -9 -6 -5
rect 112 -9 116 -5
<< metal1 >>
rect -26 170 -18 174
rect -24 158 -20 170
rect -24 132 -20 143
rect 18 142 23 152
rect 12 138 23 142
rect -24 128 -10 132
rect 18 129 23 138
rect -24 124 -20 128
rect 27 140 32 152
rect 27 136 52 140
rect 27 129 32 136
rect 48 114 52 136
rect -24 97 -20 109
rect 48 110 63 114
rect -26 93 -18 97
rect 18 86 23 98
rect 12 82 23 86
rect 18 75 23 82
rect 27 86 32 98
rect 48 86 52 110
rect 27 82 52 86
rect 27 75 32 82
rect 59 47 63 110
rect 59 43 122 47
rect -26 33 -18 37
rect 96 33 104 37
rect -24 21 -20 33
rect 98 21 102 33
rect -24 -5 -20 6
rect 18 3 23 15
rect 12 -1 23 3
rect -24 -9 -10 -5
rect 18 -8 23 -1
rect -24 -13 -20 -9
rect 27 3 32 15
rect 27 -1 52 3
rect 27 -8 32 -1
rect -24 -40 -20 -28
rect -26 -44 -18 -40
rect 18 -51 23 -39
rect 12 -55 23 -51
rect 18 -62 23 -55
rect 27 -51 32 -39
rect 48 -39 52 -1
rect 98 -5 102 6
rect 118 4 122 43
rect 140 4 145 15
rect 118 0 145 4
rect 98 -9 112 -5
rect 140 -8 145 0
rect 98 -13 102 -9
rect 149 3 154 15
rect 149 -1 174 3
rect 149 -8 154 -1
rect 170 -21 174 -1
rect 48 -43 72 -39
rect 98 -40 102 -28
rect 170 -25 182 -21
rect 48 -51 52 -43
rect 27 -55 52 -51
rect 68 -55 72 -43
rect 96 -44 104 -40
rect 140 -50 145 -39
rect 108 -54 145 -50
rect 108 -55 112 -54
rect 27 -62 32 -55
rect 68 -59 112 -55
rect 140 -62 145 -54
rect 149 -51 154 -39
rect 170 -51 174 -25
rect 149 -55 174 -51
rect 149 -62 154 -55
<< labels >>
rlabel polysilicon 81 -3 81 -3 1 S1
rlabel polysilicon -47 55 -47 55 3 S0
rlabel metal1 15 140 15 140 1 I0
rlabel metal1 15 84 15 84 1 I1
rlabel metal1 15 1 15 1 1 I2
rlabel metal1 15 -53 15 -53 1 I3
rlabel metal1 178 -23 178 -23 7 outpt
rlabel metal1 -22 172 -22 172 5 vcc
rlabel metal1 -22 95 -22 95 1 vss
rlabel metal1 -22 35 -22 35 1 vcc
rlabel metal1 -22 -42 -22 -42 1 vss
rlabel metal1 100 -42 100 -42 1 vss
rlabel metal1 100 35 100 35 1 vcc
rlabel polysilicon -2 130 -2 130 1 S0bar
<< end >>
